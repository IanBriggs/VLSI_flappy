VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  MACRO drcSignature INTEGER ;
END PROPERTYDEFINITIONS

MACRO ADDER
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN ADDER 0 0 ;
  SIZE 40.8 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN SUM
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER via ;
        RECT 39 22.5 39.6 23.1 ;
        RECT 39 2.4 39.6 3 ;
      LAYER metal2 ;
        RECT 38.7 2.1 39.9 23.4 ;
      LAYER metal1 ;
        RECT 38.7 2.1 39.9 3.3 ;
        RECT 38.7 22.2 39.9 24.9 ;
    END
  END SUM
  PIN COUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER via ;
        RECT 34.2 22.5 34.8 23.1 ;
        RECT 34.2 2.4 34.8 3 ;
      LAYER metal2 ;
        RECT 33.9 2.1 35.1 23.4 ;
      LAYER metal1 ;
        RECT 33.9 2.1 35.1 3.3 ;
        RECT 33.9 22.2 35.1 24.9 ;
    END
  END COUT
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 15.6 1.8 16.8 ;
        RECT 0.6 15.75 7.2 16.65 ;
        RECT 9 15.3 10.2 16.5 ;
        RECT 6.3 15.45 14.4 16.35 ;
        RECT 13.5 13.65 14.4 16.35 ;
        RECT 13.5 13.65 24 14.55 ;
        RECT 22.8 13.5 24 14.7 ;
    END
  END A
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3 19.5 4.2 28.2 ;
        RECT 11.7 19.5 12.9 28.2 ;
        RECT 21.3 19.5 22.5 28.2 ;
        RECT 26.1 19.5 27.3 28.2 ;
        RECT 36.3 22.5 37.5 28.2 ;
        RECT -1.2 25.8 42 28.2 ;
    END
  END vdd!
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.4 9.6 6.6 10.8 ;
        RECT 20.1 9.6 21.3 10.8 ;
        RECT 5.4 9.75 32.4 10.65 ;
        RECT 31.2 9.6 32.4 10.8 ;
    END
  END CIN
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3 -1.2 4.2 4.5 ;
        RECT 11.7 -1.2 12.9 4.5 ;
        RECT 21.3 -1.2 22.5 4.5 ;
        RECT 26.1 -1.2 27.3 4.5 ;
        RECT 36.3 -1.2 37.5 3 ;
        RECT -1.2 -1.2 42 1.2 ;
    END
  END gnd!
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 12.6 4.2 13.8 ;
        RECT 3 12.75 12 13.65 ;
        RECT 11.1 11.55 12.3 12.75 ;
        RECT 11.1 11.7 29.1 12.6 ;
        RECT 27.9 11.55 29.1 12.75 ;
    END
  END B
  OBS
    LAYER metal1 ;
      RECT 0.9 17.7 6.3 18.6 ;
      RECT 5.4 17.7 6.3 24.9 ;
      RECT 0.9 17.7 1.8 24.9 ;
      RECT 0.6 19.2 1.8 24.9 ;
      RECT 5.4 19.2 6.6 24.9 ;
      RECT 0.6 2.1 1.8 4.8 ;
      RECT 5.4 2.1 6.6 4.8 ;
      RECT 0.9 2.1 1.8 6.3 ;
      RECT 5.4 2.1 6.3 6.3 ;
      RECT 0.9 5.4 6.3 6.3 ;
      RECT 14.1 19.2 15.3 24.9 ;
      RECT 14.1 2.1 15.3 4.8 ;
      RECT 18.9 19.2 20.1 24.9 ;
      RECT 18.9 2.1 20.1 4.8 ;
      RECT 23.7 19.2 24.9 24.9 ;
      RECT 23.7 2.1 24.9 4.8 ;
      RECT 35.1 15.3 36.3 16.5 ;
      RECT 15.3 15.6 36.3 16.5 ;
      RECT 15.3 15.45 16.5 16.65 ;
      RECT 15.3 15.45 16.2 18.3 ;
      RECT 8.1 17.4 16.2 18.3 ;
      RECT 8.1 17.4 9 24.9 ;
      RECT 7.8 19.2 9 24.9 ;
      RECT 7.8 2.1 9 4.8 ;
      RECT 7.95 2.1 8.85 8.4 ;
      RECT 7.95 7.5 36.3 8.4 ;
      RECT 15.3 7.35 16.5 8.55 ;
      RECT 35.1 7.5 36.3 8.7 ;
      RECT 17.1 17.4 38.7 18.3 ;
      RECT 37.5 17.25 38.7 18.45 ;
      RECT 31.65 17.4 32.55 24.9 ;
      RECT 17.1 17.4 18 24.9 ;
      RECT 16.5 19.2 18 24.9 ;
      RECT 31.5 19.2 32.7 24.9 ;
      RECT 16.5 2.1 18 4.8 ;
      RECT 31.5 2.1 32.7 4.8 ;
      RECT 17.1 2.1 18 6.6 ;
      RECT 31.65 2.1 32.55 6.6 ;
      RECT 17.1 5.7 38.7 6.6 ;
      RECT 37.5 5.55 38.7 6.75 ;
    LAYER metal2 ;
      RECT 14.1 23.85 24.9 24.75 ;
      RECT 14.1 23.7 15.3 24.9 ;
      RECT 18.9 23.7 20.1 24.9 ;
      RECT 23.7 23.7 24.9 24.9 ;
      RECT 14.1 2.25 24.9 3.15 ;
      RECT 14.1 2.1 15.3 3.3 ;
      RECT 18.9 2.1 20.1 3.3 ;
      RECT 23.7 2.1 24.9 3.3 ;
    LAYER via ;
      RECT 14.4 24 15 24.6 ;
      RECT 14.4 2.4 15 3 ;
      RECT 19.2 24 19.8 24.6 ;
      RECT 19.2 2.4 19.8 3 ;
      RECT 24 24 24.6 24.6 ;
      RECT 24 2.4 24.6 3 ;
  END
  PROPERTY drcSignature 14016396 ;
END ADDER

MACRO AOI22
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN AOI22 0 0 ;
  SIZE 12 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER via ;
        RECT 5.7 19.5 6.3 20.1 ;
        RECT 5.7 3.9 6.3 4.5 ;
      LAYER metal2 ;
        RECT 5.4 3.6 6.6 20.4 ;
      LAYER metal1 ;
        RECT 5.4 2.1 6.6 4.8 ;
        RECT 5.4 19.2 6.6 24.9 ;
    END
  END Y
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.8 9.9 9 11.1 ;
    END
  END D
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 1.8 6.9 3 8.1 ;
        RECT 1.8 7.05 11.4 7.95 ;
        RECT 10.2 6.9 11.4 8.1 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 12.9 4.2 14.1 ;
    END
  END C
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 15.9 1.8 17.1 ;
    END
  END A
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 19.5 1.8 28.2 ;
        RECT 10.2 19.5 11.4 28.2 ;
        RECT -1.2 25.8 13.2 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 4.5 ;
        RECT 10.2 -1.2 11.4 4.5 ;
        RECT -1.2 -1.2 13.2 1.2 ;
    END
  END gnd!
  OBS
    LAYER metal1 ;
      RECT 3 2.1 4.2 4.8 ;
      RECT 3.3 17.4 8.7 18.3 ;
      RECT 7.8 17.4 8.7 24.9 ;
      RECT 3.3 17.4 4.2 24.9 ;
      RECT 3 19.2 4.2 24.9 ;
      RECT 7.8 19.2 9 24.9 ;
      RECT 7.8 2.1 9 4.8 ;
  END
  PROPERTY drcSignature 14016396 ;
END AOI22

MACRO BUFX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX4 0 0 ;
  SIZE 7.2 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3 15 4.2 28.2 ;
        RECT -1.2 25.8 8.4 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3 -1.2 4.2 6 ;
        RECT -1.2 -1.2 8.4 1.2 ;
    END
  END gnd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 9.9 1.8 11.1 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.4 2.1 6.6 24.9 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.6 2.1 2.1 3.3 ;
      RECT 1.2 2.1 2.1 7.8 ;
      RECT 1.2 6.9 4.35 7.8 ;
      RECT 3.3 9.9 4.5 11.1 ;
      RECT 3.45 6.9 4.35 14.1 ;
      RECT 1.2 13.2 4.35 14.1 ;
      RECT 1.2 13.2 2.1 24.9 ;
      RECT 0.6 22.2 2.1 24.9 ;
  END
  PROPERTY drcSignature 14016396 ;
END BUFX4

MACRO BUFX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN BUFX8 0 0 ;
  SIZE 9.6 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3 15 4.2 28.2 ;
        RECT 7.8 13.5 9 28.2 ;
        RECT -1.2 25.8 10.8 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 3 -1.2 4.2 6 ;
        RECT 7.8 -1.2 9 7.5 ;
        RECT -1.2 -1.2 10.8 1.2 ;
    END
  END gnd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 9.9 1.8 11.1 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 5.4 2.1 6.6 24.9 ;
    END
  END Y
  OBS
    LAYER metal1 ;
      RECT 0.6 2.1 2.1 3.3 ;
      RECT 1.2 2.1 2.1 7.8 ;
      RECT 1.2 6.9 4.35 7.8 ;
      RECT 3.3 9.9 4.5 11.1 ;
      RECT 3.45 6.9 4.35 14.1 ;
      RECT 1.2 13.2 4.35 14.1 ;
      RECT 1.2 13.2 2.1 24.9 ;
      RECT 0.6 22.2 2.1 24.9 ;
  END
  PROPERTY drcSignature 14016396 ;
END BUFX8

MACRO DFF
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DFF 0 0 ;
  SIZE 38.4 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER via ;
        RECT 5.7 24 6.3 24.6 ;
        RECT 5.7 22.5 6.3 23.1 ;
        RECT 5.7 21 6.3 21.6 ;
        RECT 5.7 19.5 6.3 20.1 ;
        RECT 5.7 3.9 6.3 4.5 ;
        RECT 5.7 2.4 6.3 3 ;
      LAYER metal2 ;
        RECT 5.4 2.1 6.6 24.9 ;
      LAYER metal1 ;
        RECT 5.4 2.1 6.6 4.8 ;
        RECT 5.4 19.2 6.6 24.9 ;
    END
  END D
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 3 ;
        RECT 11.7 -1.2 12.9 4.5 ;
        RECT 21.9 -1.2 23.1 4.5 ;
        RECT 26.7 -1.2 27.9 4.5 ;
        RECT 33.9 -1.2 35.1 3 ;
        RECT -1.2 -1.2 39.6 1.2 ;
    END
  END gnd!
  PIN QB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER via ;
        RECT 36.6 24 37.2 24.6 ;
        RECT 36.6 22.5 37.2 23.1 ;
        RECT 36.6 2.4 37.2 3 ;
      LAYER metal2 ;
        RECT 36.3 2.1 37.5 24.9 ;
      LAYER metal1 ;
        RECT 36.3 2.1 37.5 3.3 ;
        RECT 36.3 22.2 37.5 24.9 ;
    END
  END QB
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER via ;
        RECT 24.6 14.1 25.2 14.7 ;
        RECT 24.6 3.9 25.2 4.5 ;
        RECT 24.6 2.4 25.2 3 ;
      LAYER metal2 ;
        RECT 24.3 2.1 25.5 15 ;
      LAYER metal1 ;
        RECT 35.1 13.8 36.3 15 ;
        RECT 24.3 13.8 36.3 14.7 ;
        RECT 29.1 19.2 30.3 24.9 ;
        RECT 29.1 17.7 30 24.9 ;
        RECT 28.5 13.8 29.4 18.6 ;
        RECT 24.3 13.8 25.5 15 ;
        RECT 20.4 7.8 25.8 8.7 ;
        RECT 24.9 2.1 25.8 8.7 ;
        RECT 24.3 2.1 25.8 4.8 ;
        RECT 20.4 7.5 21.6 8.7 ;
    END
  END Q
  PIN CLRB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 14.7 9.6 33.9 10.8 ;
    END
  END CLRB
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 0.6 11.7 1.8 14.1 ;
        RECT 0.6 11.7 23.1 12.9 ;
    END
  END CLK
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 22.5 1.8 28.2 ;
        RECT 11.7 19.5 12.9 28.2 ;
        RECT 16.5 22.5 17.7 28.2 ;
        RECT 25.2 19.5 26.4 28.2 ;
        RECT 33.9 22.5 35.1 28.2 ;
        RECT -1.2 25.8 39.6 28.2 ;
    END
  END vdd!
  OBS
    LAYER metal1 ;
      RECT 3 2.1 4.2 3.3 ;
      RECT 3.3 2.1 4.2 8.7 ;
      RECT 3.3 7.5 4.5 8.7 ;
      RECT 12.6 17.4 13.8 18.6 ;
      RECT 8.1 17.7 13.8 18.6 ;
      RECT 8.1 17.7 9 24.9 ;
      RECT 7.8 19.2 9 24.9 ;
      RECT 7.8 2.1 9 4.8 ;
      RECT 8.1 2.1 9 6.45 ;
      RECT 8.1 5.55 13.8 6.45 ;
      RECT 12.6 5.55 13.8 6.75 ;
      RECT 15.6 2.1 16.8 3.3 ;
      RECT 10.2 7.5 11.4 8.7 ;
      RECT 15.75 2.1 16.65 8.7 ;
      RECT 10.2 7.8 16.65 8.7 ;
      RECT 10.2 15.6 18.9 16.5 ;
      RECT 10.2 15.6 11.4 16.8 ;
      RECT 18 15.6 18.9 20.25 ;
      RECT 14.4 19.35 20.1 20.25 ;
      RECT 14.4 19.35 15.3 24.9 ;
      RECT 14.1 22.2 15.3 24.9 ;
      RECT 18.9 19.2 20.1 24.9 ;
      RECT 3.3 13.8 21 14.7 ;
      RECT 3.3 13.8 4.5 15 ;
      RECT 8.1 13.8 9.3 15 ;
      RECT 19.8 13.8 21 15 ;
      RECT 3.3 13.8 4.2 24.9 ;
      RECT 3 22.2 4.2 24.9 ;
      RECT 18 2.1 19.2 4.8 ;
      RECT 18.15 2.1 19.05 6.6 ;
      RECT 18.15 5.7 24 6.6 ;
      RECT 22.8 5.7 24 6.9 ;
      RECT 26.4 15.6 27.6 16.8 ;
      RECT 21.45 15.9 27.6 16.8 ;
      RECT 21.45 15.9 22.35 24.9 ;
      RECT 21.3 19.2 22.5 24.9 ;
      RECT 29.1 2.1 30.3 3.3 ;
      RECT 29.1 2.4 31.35 3.3 ;
      RECT 30.45 2.4 31.35 8.7 ;
      RECT 30.3 7.5 31.5 8.7 ;
      RECT 30.3 15.6 31.5 16.8 ;
      RECT 30.3 15.9 32.55 16.8 ;
      RECT 31.65 15.9 32.55 24.9 ;
      RECT 31.5 22.2 32.7 24.9 ;
  END
  PROPERTY drcSignature 14016396 ;
END DFF

MACRO FILLER
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN FILLER 0 0 ;
  SIZE 2.4 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.05 -1.2 1.95 1.8 ;
        RECT -1.2 -1.2 3.6 1.2 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.05 25.2 1.95 28.2 ;
        RECT -1.2 25.8 3.6 28.2 ;
    END
  END vdd!
  PROPERTY drcSignature 14016396 ;
END FILLER

MACRO INVX1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX1 0 0 ;
  SIZE 4.8 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 22.5 1.8 28.2 ;
        RECT -1.2 25.8 6 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 3 ;
        RECT -1.2 -1.2 6 1.2 ;
    END
  END gnd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.9 9.9 2.1 11.1 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 2.1 4.2 24.9 ;
    END
  END Y
  PROPERTY drcSignature 14016396 ;
END INVX1

MACRO INVX4
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX4 0 0 ;
  SIZE 4.8 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 13.5 1.8 28.2 ;
        RECT -1.2 25.8 6 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 7.5 ;
        RECT -1.2 -1.2 6 1.2 ;
    END
  END gnd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.9 9.9 2.1 11.1 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 2.1 4.2 24.9 ;
    END
  END Y
  PROPERTY drcSignature 14016396 ;
END INVX4

MACRO INVX8
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN INVX8 0 0 ;
  SIZE 7.2 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 13.5 1.8 28.2 ;
        RECT 5.4 13.5 6.6 28.2 ;
        RECT -1.2 25.8 8.4 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 7.5 ;
        RECT 5.4 -1.2 6.6 7.5 ;
        RECT -1.2 -1.2 8.4 1.2 ;
    END
  END gnd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.9 9.9 2.1 11.1 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 2.1 4.2 24.9 ;
    END
  END Y
  PROPERTY drcSignature 14016396 ;
END INVX8

MACRO MUX2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN MUX2X1 0 0 ;
  SIZE 12 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 4.2 -1.2 5.7 1.8 ;
        RECT 4.5 -1.2 5.7 4.5 ;
        RECT -1.2 -1.2 13.2 1.2 ;
    END
  END gnd!
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 4.5 19.5 5.7 28.2 ;
        RECT 4.2 25.2 5.7 28.2 ;
        RECT -1.2 25.8 13.2 28.2 ;
    END
  END vdd!
  PIN D0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.45 12.9 1.65 14.1 ;
    END
  END D0
  PIN D1
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.95 7.2 9.15 8.4 ;
    END
  END D1
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.3 15.6 4.5 16.8 ;
        RECT 5.85 9.9 6.75 16.5 ;
        RECT 3.3 15.6 6.75 16.5 ;
        RECT 5.7 9.9 6.9 11.1 ;
    END
  END S
  PIN SB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.3 9.9 4.5 11.1 ;
    END
  END SB
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 2.1 1.8 4.8 ;
        RECT 0.9 2.1 1.8 6.3 ;
        RECT 0.9 17.7 1.8 24.9 ;
        RECT 0.6 19.2 1.8 24.9 ;
        RECT 0.9 17.7 9.3 18.6 ;
        RECT 8.4 2.1 9.3 6.3 ;
        RECT 0.9 5.4 9.3 6.3 ;
        RECT 8.4 17.7 9.3 24.9 ;
        RECT 8.4 2.1 9.6 4.8 ;
        RECT 8.4 19.2 9.6 24.9 ;
        RECT 8.4 3.6 11.4 4.8 ;
        RECT 10.2 3.6 11.4 20.4 ;
        RECT 8.4 19.2 11.4 20.4 ;
    END
  END Y
  PROPERTY drcSignature 14016396 ;
END MUX2X1

MACRO NAND2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X1 0 0 ;
  SIZE 7.2 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 20.4 4.2 24.9 ;
        RECT 4.8 2.1 6.6 4.8 ;
        RECT 5.4 2.1 6.6 21.6 ;
        RECT 3 20.4 6.6 21.6 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 9.9 4.2 11.1 ;
    END
  END B
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.9 -1.2 2.1 4.5 ;
        RECT -1.2 -1.2 8.4 1.2 ;
    END
  END gnd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 12.9 1.8 14.1 ;
    END
  END A
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 22.5 1.8 28.2 ;
        RECT 5.4 22.5 6.6 28.2 ;
        RECT -1.2 25.8 8.4 28.2 ;
    END
  END vdd!
  PROPERTY drcSignature 14016396 ;
END NAND2X1

MACRO NAND2X2
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NAND2X2 0 0 ;
  SIZE 7.2 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 17.4 4.2 24.9 ;
        RECT 4.8 2.1 6.6 7.8 ;
        RECT 5.4 2.1 6.6 18.6 ;
        RECT 3 17.4 6.6 18.6 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 9.9 4.2 11.1 ;
    END
  END B
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.9 -1.2 2.1 7.5 ;
        RECT -1.2 -1.2 8.4 1.2 ;
    END
  END gnd!
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 12.9 1.8 14.1 ;
    END
  END A
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 19.5 1.8 28.2 ;
        RECT 5.4 19.5 6.6 28.2 ;
        RECT -1.2 25.8 8.4 28.2 ;
    END
  END vdd!
  PROPERTY drcSignature 14016396 ;
END NAND2X2

MACRO NOR2X1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN NOR2X1 0 0 ;
  SIZE 7.2 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 2.1 4.2 5.1 ;
        RECT 3 3.9 6.6 5.1 ;
        RECT 5.4 3.9 6.6 24.9 ;
        RECT 4.8 19.2 6.6 24.9 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 9.9 4.2 11.1 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 12.9 1.8 14.1 ;
    END
  END A
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.9 19.5 2.1 28.2 ;
        RECT -1.2 25.8 8.4 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 3 ;
        RECT 5.4 -1.2 6.6 3 ;
        RECT -1.2 -1.2 8.4 1.2 ;
    END
  END gnd!
  PROPERTY drcSignature 14016396 ;
END NOR2X1

MACRO OAI22
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN OAI22 0 0 ;
  SIZE 12 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER via ;
        RECT 5.7 19.5 6.3 20.1 ;
        RECT 5.7 3.9 6.3 4.5 ;
      LAYER metal2 ;
        RECT 5.4 3.6 6.6 20.4 ;
      LAYER metal1 ;
        RECT 5.4 2.1 6.6 4.8 ;
        RECT 5.4 19.2 6.6 24.9 ;
    END
  END Y
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 9.9 4.2 11.1 ;
        RECT 9 8.1 9.9 10.8 ;
        RECT 3 9.9 9.9 10.8 ;
        RECT 9 8.1 10.2 9.3 ;
    END
  END C
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 10.2 15.9 11.4 17.1 ;
    END
  END B
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 6.9 1.8 8.1 ;
    END
  END D
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 7.8 12.9 9 14.1 ;
    END
  END A
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 19.5 1.8 28.2 ;
        RECT 10.2 19.5 11.4 28.2 ;
        RECT -1.2 25.8 13.2 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 4.5 ;
        RECT 10.2 -1.2 11.4 4.5 ;
        RECT -1.2 -1.2 13.2 1.2 ;
    END
  END gnd!
  OBS
    LAYER metal1 ;
      RECT 3 19.2 4.2 24.9 ;
      RECT 7.8 19.2 9 24.9 ;
      RECT 3 2.1 4.2 4.8 ;
      RECT 7.8 2.1 9 4.8 ;
      RECT 3.3 2.1 4.2 6.6 ;
      RECT 7.8 2.1 8.7 6.6 ;
      RECT 3.3 5.7 8.7 6.6 ;
  END
  PROPERTY drcSignature 14016396 ;
END OAI22

MACRO TIEHI
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIEHI 0 0 ;
  SIZE 4.8 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 19.2 4.2 24.9 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 19.5 1.8 28.2 ;
        RECT -1.2 25.8 6 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 4.5 ;
        RECT -1.2 -1.2 6 1.2 ;
    END
  END gnd!
  OBS
    LAYER metal1 ;
      RECT 3 2.1 4.2 6.9 ;
      RECT 1.8 5.7 4.2 6.9 ;
  END
  PROPERTY drcSignature 14016396 ;
END TIEHI

MACRO TIELO
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN TIELO 0 0 ;
  SIZE 4.8 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 2.1 4.2 4.8 ;
    END
  END Y
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 19.5 1.8 28.2 ;
        RECT -1.2 25.8 6 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 4.5 ;
        RECT -1.2 -1.2 6 1.2 ;
    END
  END gnd!
  OBS
    LAYER metal1 ;
      RECT 1.8 17.1 4.2 18.3 ;
      RECT 3 17.1 4.2 24.9 ;
  END
  PROPERTY drcSignature 14016396 ;
END TIELO

MACRO XOR
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN XOR 0 0 ;
  SIZE 19.2 BY 27 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 11.7 2.1 14.1 4.8 ;
        RECT 11.7 17.4 12.9 24.9 ;
        RECT 12.9 2.1 14.1 6.6 ;
        RECT 12.9 5.4 16.8 6.6 ;
        RECT 15.6 5.4 16.8 18.6 ;
        RECT 11.7 17.4 16.8 18.6 ;
    END
  END Y
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3 9.9 4.2 11.1 ;
        RECT 3 10.05 14.1 10.95 ;
        RECT 12.9 10.05 14.1 12.15 ;
    END
  END B
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.6 12.9 1.8 14.1 ;
        RECT 0.6 13.05 10.8 13.95 ;
        RECT 9.6 12.9 10.8 14.1 ;
    END
  END A
  PIN vdd!
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 22.5 1.8 28.2 ;
        RECT 7.8 19.5 9 28.2 ;
        RECT 15.6 19.5 16.8 28.2 ;
        RECT -1.2 25.8 20.4 28.2 ;
    END
  END vdd!
  PIN gnd!
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 0.6 -1.2 1.8 3 ;
        RECT 7.8 -1.2 9 4.5 ;
        RECT 15.6 -1.2 16.8 4.5 ;
        RECT -1.2 -1.2 20.4 1.2 ;
    END
  END gnd!
  OBS
    LAYER metal1 ;
      RECT 4.8 15.3 6 16.5 ;
      RECT 3.15 15.6 6 16.5 ;
      RECT 3.15 15.6 4.05 24.9 ;
      RECT 3 22.2 4.2 24.9 ;
      RECT 3 2.1 4.2 3.3 ;
      RECT 3.15 2.1 4.05 8.7 ;
      RECT 3.15 7.8 6 8.7 ;
      RECT 4.8 7.8 6 9 ;
      RECT 5.4 2.1 6.6 3.3 ;
      RECT 5.7 2.1 6.6 6.9 ;
      RECT 5.7 6 12 6.9 ;
      RECT 10.8 6 12 7.5 ;
      RECT 12.6 15.3 13.8 16.5 ;
      RECT 7.95 15.6 13.8 16.5 ;
      RECT 7.95 15.6 8.85 18.3 ;
      RECT 5.55 17.4 8.85 18.3 ;
      RECT 5.55 17.4 6.45 24.9 ;
      RECT 5.4 22.2 6.6 24.9 ;
  END
  PROPERTY drcSignature 14016396 ;
END XOR

END LIBRARY
